LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
  
PACKAGE type_pkg IS  
  --TYPE STATE IS (INIT, LOAD, RE_LOAD, SHIFT, DONE);
  SUBTYPE SLV_8 IS STD_LOGIC_VECTOR(7 DOWNTO 0); 
  SUBTYPE STATE_TYPE IS STD_LOGIC_VECTOR(127 DOWNTO 0); 
  SUBTYPE SLV_128 IS STD_LOGIC_VECTOR(127 DOWNTO 0); 
  SUBTYPE SLV_32 IS STD_LOGIC_VECTOR(31 DOWNTO 0); 
  SUBTYPE ROUND_TYPE IS INTEGER RANGE 0 TO 16;
  TYPE STATE_ARRAY IS ARRAY (15 DOWNTO 0) OF SLV_8;
  TYPE STATE_ARRAY2 IS ARRAY (10 DOWNTO 0) OF STATE_ARRAY;
  TYPE COLUMN_STATE_ARRAY IS ARRAY (3 DOWNTO 0) OF SLV_8;
END PACKAGE type_pkg; 
