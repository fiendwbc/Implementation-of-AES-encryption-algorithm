LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE work.ALL;
USE work.type_pkg.ALL;

ENTITY multiplier_substitute IS
    PORT(a, b: IN SLV_8; c: OUT SLV_8);
END multiplier_substitute;
  
ARCHITECTURE rtl OF multiplier_substitute IS
  COMPONENT sbox_lookup
      PORT(a: IN SLV_8; b: OUT SLV_8);
  END COMPONENT;
 -- SIGNAL cWord: SLV_8;
 -- SIGNAL b: SLV_8;
 -- SIGNAL cIndex: INTEGER :=0;
 -- SIGNAL t: STATE_ARRAY;
BEGIN
  find:PROCESS(a, b)
  BEGIN
		CASE a IS
		WHEN x"09" =>
			CASE b IS
				WHEN x"00" => c <= x"00"; 
				WHEN x"01" => c <= x"09"; 
				WHEN x"02" => c <= x"12"; 
				WHEN x"03" => c <= x"1b"; 
				WHEN x"04" => c <= x"24"; 
				WHEN x"05" => c <= x"2d"; 
				WHEN x"06" => c <= x"36"; 
				WHEN x"07" => c <= x"3f"; 
				WHEN x"08" => c <= x"48"; 
				WHEN x"09" => c <= x"41"; 
				WHEN x"0a" => c <= x"5a"; 
				WHEN x"0b" => c <= x"53"; 
				WHEN x"0c" => c <= x"6c"; 
				WHEN x"0d" => c <= x"65"; 
				WHEN x"0e" => c <= x"7e"; 
				WHEN x"0f" => c <= x"77";  
				WHEN x"10" => c <= x"90"; 
				WHEN x"11" => c <= x"99"; 
				WHEN x"12" => c <= x"82"; 
				WHEN x"13" => c <= x"8b"; 
				WHEN x"14" => c <= x"b4"; 
				WHEN x"15" => c <= x"bd"; 
				WHEN x"16" => c <= x"a6"; 
				WHEN x"17" => c <= x"af"; 
				WHEN x"18" => c <= x"d8"; 
				WHEN x"19" => c <= x"d1"; 
				WHEN x"1a" => c <= x"ca"; 
				WHEN x"1b" => c <= x"c3"; 
				WHEN x"1c" => c <= x"fc"; 
				WHEN x"1d" => c <= x"f5"; 
				WHEN x"1e" => c <= x"ee"; 
				WHEN x"1f" => c <= x"e7";
				WHEN x"20" => c <= x"3b";
				WHEN x"21" => c <= x"32"; 
				WHEN x"22" => c <= x"29"; 
				WHEN x"23" => c <= x"20"; 
				WHEN x"24" => c <= x"1f"; 
				WHEN x"25" => c <= x"16"; 
				WHEN x"26" => c <= x"0d"; 
				WHEN x"27" => c <= x"04"; 
				WHEN x"28" => c <= x"73"; 
				WHEN x"29" => c <= x"7a"; 
				WHEN x"2a" => c <= x"61"; 
				WHEN x"2b" => c <= x"68"; 
				WHEN x"2c" => c <= x"57"; 
				WHEN x"2d" => c <= x"5e"; 
				WHEN x"2e" => c <= x"45"; 
				WHEN x"2f" => c <= x"4c";  
				WHEN x"30" => c <= x"ab"; 
				WHEN x"31" => c <= x"a2"; 
				WHEN x"32" => c <= x"b9"; 
				WHEN x"33" => c <= x"b0"; 
				WHEN x"34" => c <= x"8f"; 
				WHEN x"35" => c <= x"86"; 
				WHEN x"36" => c <= x"9d"; 
				WHEN x"37" => c <= x"94"; 
				WHEN x"38" => c <= x"e3"; 
				WHEN x"39" => c <= x"ea"; 
				WHEN x"3a" => c <= x"f1"; 
				WHEN x"3b" => c <= x"f8"; 
				WHEN x"3c" => c <= x"c7"; 
				WHEN x"3d" => c <= x"ce"; 
				WHEN x"3e" => c <= x"d5"; 
				WHEN x"3f" => c <= x"dc";
				WHEN x"40" => c <= x"76"; 
				WHEN x"41" => c <= x"7f"; 
				WHEN x"42" => c <= x"64"; 
				WHEN x"43" => c <= x"6d"; 
				WHEN x"44" => c <= x"52"; 
				WHEN x"45" => c <= x"5b"; 
				WHEN x"46" => c <= x"40"; 
				WHEN x"47" => c <= x"49"; 
				WHEN x"48" => c <= x"3e"; 
				WHEN x"49" => c <= x"37"; 
				WHEN x"4a" => c <= x"2c"; 
				WHEN x"4b" => c <= x"25"; 
				WHEN x"4c" => c <= x"1a"; 
				WHEN x"4d" => c <= x"13"; 
				WHEN x"4e" => c <= x"08"; 
				WHEN x"4f" => c <= x"01";  
				WHEN x"50" => c <= x"e6";
				WHEN x"51" => c <= x"ef";
				WHEN x"52" => c <= x"f4";
				WHEN x"53" => c <= x"fd";
				WHEN x"54" => c <= x"c2";
				WHEN x"55" => c <= x"cb";
				WHEN x"56" => c <= x"d0";
				WHEN x"57" => c <= x"d9";
				WHEN x"58" => c <= x"ae";
				WHEN x"59" => c <= x"a7";
				WHEN x"5a" => c <= x"bc";
				WHEN x"5b" => c <= x"b5";
				WHEN x"5c" => c <= x"8a";
				WHEN x"5d" => c <= x"83";
				WHEN x"5e" => c <= x"98";
				WHEN x"5f" => c <= x"91"; 
				WHEN x"60" => c <= x"4d";
				WHEN x"61" => c <= x"44";
				WHEN x"62" => c <= x"5f";
				WHEN x"63" => c <= x"56";
				WHEN x"64" => c <= x"69";
				WHEN x"65" => c <= x"60";
				WHEN x"66" => c <= x"7b";
				WHEN x"67" => c <= x"72";
				WHEN x"68" => c <= x"05";
				WHEN x"69" => c <= x"0c";
				WHEN x"6a" => c <= x"17";
				WHEN x"6b" => c <= x"1e";
				WHEN x"6c" => c <= x"21";
				WHEN x"6d" => c <= x"28";
				WHEN x"6e" => c <= x"33";
				WHEN x"6f" => c <= x"3a";  
				WHEN x"70" => c <= x"dd";
				WHEN x"71" => c <= x"d4";
				WHEN x"72" => c <= x"cf";
				WHEN x"73" => c <= x"c6";
				WHEN x"74" => c <= x"f9";
				WHEN x"75" => c <= x"f0";
				WHEN x"76" => c <= x"eb";
				WHEN x"77" => c <= x"e2";
				WHEN x"78" => c <= x"95";
				WHEN x"79" => c <= x"9c";
				WHEN x"7a" => c <= x"87";
				WHEN x"7b" => c <= x"8e";
				WHEN x"7c" => c <= x"b1";
				WHEN x"7d" => c <= x"b8";
				WHEN x"7e" => c <= x"a3";
				WHEN x"7f" => c <= x"aa"; 
				WHEN x"80" => c <= x"ec";
				WHEN x"81" => c <= x"e5";
				WHEN x"82" => c <= x"fe";
				WHEN x"83" => c <= x"f7";
				WHEN x"84" => c <= x"c8";
				WHEN x"85" => c <= x"c1";
				WHEN x"86" => c <= x"da";
				WHEN x"87" => c <= x"d3";
				WHEN x"88" => c <= x"a4";
				WHEN x"89" => c <= x"ad";
				WHEN x"8a" => c <= x"b6";
				WHEN x"8b" => c <= x"bf";
				WHEN x"8c" => c <= x"80";
				WHEN x"8d" => c <= x"89";
				WHEN x"8e" => c <= x"92";
				WHEN x"8f" => c <= x"9b";  
				WHEN x"90" => c <= x"7c";
				WHEN x"91" => c <= x"75";
				WHEN x"92" => c <= x"6e";
				WHEN x"93" => c <= x"67";
				WHEN x"94" => c <= x"58";
				WHEN x"95" => c <= x"51";
				WHEN x"96" => c <= x"4a";
				WHEN x"97" => c <= x"43";
				WHEN x"98" => c <= x"34";
				WHEN x"99" => c <= x"3d";
				WHEN x"9a" => c <= x"26";
				WHEN x"9b" => c <= x"2f";
				WHEN x"9c" => c <= x"10";
				WHEN x"9d" => c <= x"19";
				WHEN x"9e" => c <= x"02";
				WHEN x"9f" => c <= x"0b"; 
				WHEN x"a0" => c <= x"d7";
				WHEN x"a1" => c <= x"de";
				WHEN x"a2" => c <= x"c5";
				WHEN x"a3" => c <= x"cc";
				WHEN x"a4" => c <= x"f3";
				WHEN x"a5" => c <= x"fa";
				WHEN x"a6" => c <= x"e1";
				WHEN x"a7" => c <= x"e8";
				WHEN x"a8" => c <= x"9f";
				WHEN x"a9" => c <= x"96";
				WHEN x"aa" => c <= x"8d";
				WHEN x"ab" => c <= x"84";
				WHEN x"ac" => c <= x"bb";
				WHEN x"ad" => c <= x"b2";
				WHEN x"ae" => c <= x"a9";
				WHEN x"af" => c <= x"a0";  
				WHEN x"b0" => c <= x"47";
				WHEN x"b1" => c <= x"4e";
				WHEN x"b2" => c <= x"55";
				WHEN x"b3" => c <= x"5c";
				WHEN x"b4" => c <= x"63";
				WHEN x"b5" => c <= x"6a";
				WHEN x"b6" => c <= x"71";
				WHEN x"b7" => c <= x"78";
				WHEN x"b8" => c <= x"0f";
				WHEN x"b9" => c <= x"06";
				WHEN x"ba" => c <= x"1d";
				WHEN x"bb" => c <= x"14";
				WHEN x"bc" => c <= x"2b";
				WHEN x"bd" => c <= x"22";
				WHEN x"be" => c <= x"39";
				WHEN x"bf" => c <= x"30";
				WHEN x"c0" => c <= x"9a";
				WHEN x"c1" => c <= x"93";
				WHEN x"c2" => c <= x"88";
				WHEN x"c3" => c <= x"81";
				WHEN x"c4" => c <= x"be";
				WHEN x"c5" => c <= x"b7";
				WHEN x"c6" => c <= x"ac";
				WHEN x"c7" => c <= x"a5";
				WHEN x"c8" => c <= x"d2";
				WHEN x"c9" => c <= x"db";
				WHEN x"ca" => c <= x"c0";
				WHEN x"cb" => c <= x"c9";
				WHEN x"cc" => c <= x"f6";
				WHEN x"cd" => c <= x"ff";
				WHEN x"ce" => c <= x"e4";
				WHEN x"cf" => c <= x"ed";  
				WHEN x"d0" => c <= x"0a";
				WHEN x"d1" => c <= x"03";
				WHEN x"d2" => c <= x"18";
				WHEN x"d3" => c <= x"11";
				WHEN x"d4" => c <= x"2e";
				WHEN x"d5" => c <= x"27";
				WHEN x"d6" => c <= x"3c";
				WHEN x"d7" => c <= x"35";
				WHEN x"d8" => c <= x"42";
				WHEN x"d9" => c <= x"4b";
				WHEN x"da" => c <= x"50";
				WHEN x"db" => c <= x"59";
				WHEN x"dc" => c <= x"66";
				WHEN x"dd" => c <= x"6f";
				WHEN x"de" => c <= x"74";
				WHEN x"df" => c <= x"7d"; 
				WHEN x"e0" => c <= x"a1";
				WHEN x"e1" => c <= x"a8";
				WHEN x"e2" => c <= x"b3";
				WHEN x"e3" => c <= x"ba";
				WHEN x"e4" => c <= x"85";
				WHEN x"e5" => c <= x"8c";
				WHEN x"e6" => c <= x"97";
				WHEN x"e7" => c <= x"9e";
				WHEN x"e8" => c <= x"e9";
				WHEN x"e9" => c <= x"e0";
				WHEN x"ea" => c <= x"fb";
				WHEN x"eb" => c <= x"f2";
				WHEN x"ec" => c <= x"cd";
				WHEN x"ed" => c <= x"c4";
				WHEN x"ee" => c <= x"df";
				WHEN x"ef" => c <= x"d6";  
				WHEN x"f0" => c <= x"31";
				WHEN x"f1" => c <= x"38";
				WHEN x"f2" => c <= x"23";
				WHEN x"f3" => c <= x"2a";
				WHEN x"f4" => c <= x"15";
				WHEN x"f5" => c <= x"1c";
				WHEN x"f6" => c <= x"07";
				WHEN x"f7" => c <= x"0e";
				WHEN x"f8" => c <= x"79";
				WHEN x"f9" => c <= x"70";
				WHEN x"fa" => c <= x"6b";
				WHEN x"fb" => c <= x"62";
				WHEN x"fc" => c <= x"5d";
				WHEN x"fd" => c <= x"54";
				WHEN x"fe" => c <= x"4f";
				WHEN x"ff" => c <= x"46";  
				WHEN others => null;  
			END CASE; 
		WHEN x"11" =>
			CASE b IS
				WHEN x"00" => c <= x"00"; 
				WHEN x"01" => c <= x"0b"; 
				WHEN x"02" => c <= x"16"; 
				WHEN x"03" => c <= x"1d"; 
				WHEN x"04" => c <= x"2c"; 
				WHEN x"05" => c <= x"27"; 
				WHEN x"06" => c <= x"3a"; 
				WHEN x"07" => c <= x"31"; 
				WHEN x"08" => c <= x"58"; 
				WHEN x"09" => c <= x"53"; 
				WHEN x"0a" => c <= x"4e"; 
				WHEN x"0b" => c <= x"45"; 
				WHEN x"0c" => c <= x"74"; 
				WHEN x"0d" => c <= x"7f"; 
				WHEN x"0e" => c <= x"62"; 
				WHEN x"0f" => c <= x"69";  
				WHEN x"10" => c <= x"b0"; 
				WHEN x"11" => c <= x"bb"; 
				WHEN x"12" => c <= x"a6"; 
				WHEN x"13" => c <= x"ad"; 
				WHEN x"14" => c <= x"9c"; 
				WHEN x"15" => c <= x"97"; 
				WHEN x"16" => c <= x"8a"; 
				WHEN x"17" => c <= x"81"; 
				WHEN x"18" => c <= x"e8"; 
				WHEN x"19" => c <= x"e3"; 
				WHEN x"1a" => c <= x"fe"; 
				WHEN x"1b" => c <= x"f5"; 
				WHEN x"1c" => c <= x"c4"; 
				WHEN x"1d" => c <= x"cf"; 
				WHEN x"1e" => c <= x"d2"; 
				WHEN x"1f" => c <= x"d9";
				WHEN x"20" => c <= x"7b";
				WHEN x"21" => c <= x"70"; 
				WHEN x"22" => c <= x"6d"; 
				WHEN x"23" => c <= x"66"; 
				WHEN x"24" => c <= x"57"; 
				WHEN x"25" => c <= x"5c"; 
				WHEN x"26" => c <= x"41"; 
				WHEN x"27" => c <= x"4a"; 
				WHEN x"28" => c <= x"23"; 
				WHEN x"29" => c <= x"28"; 
				WHEN x"2a" => c <= x"35"; 
				WHEN x"2b" => c <= x"3e"; 
				WHEN x"2c" => c <= x"0f"; 
				WHEN x"2d" => c <= x"04"; 
				WHEN x"2e" => c <= x"19"; 
				WHEN x"2f" => c <= x"12";  
				WHEN x"30" => c <= x"cb"; 
				WHEN x"31" => c <= x"c0"; 
				WHEN x"32" => c <= x"dd"; 
				WHEN x"33" => c <= x"d6"; 
				WHEN x"34" => c <= x"e7"; 
				WHEN x"35" => c <= x"ec"; 
				WHEN x"36" => c <= x"f1"; 
				WHEN x"37" => c <= x"fa"; 
				WHEN x"38" => c <= x"93"; 
				WHEN x"39" => c <= x"98"; 
				WHEN x"3a" => c <= x"85"; 
				WHEN x"3b" => c <= x"8e"; 
				WHEN x"3c" => c <= x"bf"; 
				WHEN x"3d" => c <= x"b4"; 
				WHEN x"3e" => c <= x"a9"; 
				WHEN x"3f" => c <= x"a2";
				WHEN x"40" => c <= x"f6"; 
				WHEN x"41" => c <= x"fd"; 
				WHEN x"42" => c <= x"e0"; 
				WHEN x"43" => c <= x"eb"; 
				WHEN x"44" => c <= x"da"; 
				WHEN x"45" => c <= x"d1"; 
				WHEN x"46" => c <= x"cc"; 
				WHEN x"47" => c <= x"c7"; 
				WHEN x"48" => c <= x"ae"; 
				WHEN x"49" => c <= x"a5"; 
				WHEN x"4a" => c <= x"b8"; 
				WHEN x"4b" => c <= x"b3"; 
				WHEN x"4c" => c <= x"82"; 
				WHEN x"4d" => c <= x"89"; 
				WHEN x"4e" => c <= x"94"; 
				WHEN x"4f" => c <= x"9f";  
				WHEN x"50" => c <= x"46";
				WHEN x"51" => c <= x"4d";
				WHEN x"52" => c <= x"50";
				WHEN x"53" => c <= x"5b";
				WHEN x"54" => c <= x"6a";
				WHEN x"55" => c <= x"61";
				WHEN x"56" => c <= x"7c";
				WHEN x"57" => c <= x"77";
				WHEN x"58" => c <= x"1e";
				WHEN x"59" => c <= x"15";
				WHEN x"5a" => c <= x"08";
				WHEN x"5b" => c <= x"03";
				WHEN x"5c" => c <= x"32";
				WHEN x"5d" => c <= x"39";
				WHEN x"5e" => c <= x"24";
				WHEN x"5f" => c <= x"2f"; 
				WHEN x"60" => c <= x"8d";
				WHEN x"61" => c <= x"86";
				WHEN x"62" => c <= x"9b";
				WHEN x"63" => c <= x"90";
				WHEN x"64" => c <= x"a1";
				WHEN x"65" => c <= x"aa";
				WHEN x"66" => c <= x"b7";
				WHEN x"67" => c <= x"bc";
				WHEN x"68" => c <= x"d5";
				WHEN x"69" => c <= x"de";
				WHEN x"6a" => c <= x"c3";
				WHEN x"6b" => c <= x"c8";
				WHEN x"6c" => c <= x"f9";
				WHEN x"6d" => c <= x"f2";
				WHEN x"6e" => c <= x"ef";
				WHEN x"6f" => c <= x"e4";  
				WHEN x"70" => c <= x"3d";
				WHEN x"71" => c <= x"36";
				WHEN x"72" => c <= x"2b";
				WHEN x"73" => c <= x"20";
				WHEN x"74" => c <= x"11";
				WHEN x"75" => c <= x"1a";
				WHEN x"76" => c <= x"07";
				WHEN x"77" => c <= x"0c";
				WHEN x"78" => c <= x"65";
				WHEN x"79" => c <= x"6e";
				WHEN x"7a" => c <= x"73";
				WHEN x"7b" => c <= x"78";
				WHEN x"7c" => c <= x"49";
				WHEN x"7d" => c <= x"42";
				WHEN x"7e" => c <= x"5f";
				WHEN x"7f" => c <= x"54"; 
				WHEN x"80" => c <= x"f7";
				WHEN x"81" => c <= x"fc";
				WHEN x"82" => c <= x"e1";
				WHEN x"83" => c <= x"ea";
				WHEN x"84" => c <= x"db";
				WHEN x"85" => c <= x"d0";
				WHEN x"86" => c <= x"cd";
				WHEN x"87" => c <= x"c6";
				WHEN x"88" => c <= x"af";
				WHEN x"89" => c <= x"a4";
				WHEN x"8a" => c <= x"b9";
				WHEN x"8b" => c <= x"b2";
				WHEN x"8c" => c <= x"83";
				WHEN x"8d" => c <= x"88";
				WHEN x"8e" => c <= x"95";
				WHEN x"8f" => c <= x"9e";  
				WHEN x"90" => c <= x"47";
				WHEN x"91" => c <= x"4c";
				WHEN x"92" => c <= x"51";
				WHEN x"93" => c <= x"5a";
				WHEN x"94" => c <= x"6b";
				WHEN x"95" => c <= x"60";
				WHEN x"96" => c <= x"7d";
				WHEN x"97" => c <= x"76";
				WHEN x"98" => c <= x"1f";
				WHEN x"99" => c <= x"14";
				WHEN x"9a" => c <= x"09";
				WHEN x"9b" => c <= x"02";
				WHEN x"9c" => c <= x"33";
				WHEN x"9d" => c <= x"38";
				WHEN x"9e" => c <= x"25";
				WHEN x"9f" => c <= x"2e"; 
				WHEN x"a0" => c <= x"8c";
				WHEN x"a1" => c <= x"87";
				WHEN x"a2" => c <= x"9a";
				WHEN x"a3" => c <= x"91";
				WHEN x"a4" => c <= x"a0";
				WHEN x"a5" => c <= x"ab";
				WHEN x"a6" => c <= x"b6";
				WHEN x"a7" => c <= x"bd";
				WHEN x"a8" => c <= x"d4";
				WHEN x"a9" => c <= x"df";
				WHEN x"aa" => c <= x"c2";
				WHEN x"ab" => c <= x"c9";
				WHEN x"ac" => c <= x"f8";
				WHEN x"ad" => c <= x"f3";
				WHEN x"ae" => c <= x"ee";
				WHEN x"af" => c <= x"e5";  
				WHEN x"b0" => c <= x"3c";
				WHEN x"b1" => c <= x"37";
				WHEN x"b2" => c <= x"2a";
				WHEN x"b3" => c <= x"21";
				WHEN x"b4" => c <= x"10";
				WHEN x"b5" => c <= x"1b";
				WHEN x"b6" => c <= x"06";
				WHEN x"b7" => c <= x"0d";
				WHEN x"b8" => c <= x"64";
				WHEN x"b9" => c <= x"6f";
				WHEN x"ba" => c <= x"72";
				WHEN x"bb" => c <= x"79";
				WHEN x"bc" => c <= x"48";
				WHEN x"bd" => c <= x"43";
				WHEN x"be" => c <= x"5e";
				WHEN x"bf" => c <= x"55";
				WHEN x"c0" => c <= x"01";
				WHEN x"c1" => c <= x"0a";
				WHEN x"c2" => c <= x"17";
				WHEN x"c3" => c <= x"1c";
				WHEN x"c4" => c <= x"2d";
				WHEN x"c5" => c <= x"26";
				WHEN x"c6" => c <= x"3b";
				WHEN x"c7" => c <= x"30";
				WHEN x"c8" => c <= x"59";
				WHEN x"c9" => c <= x"52";
				WHEN x"ca" => c <= x"4f";
				WHEN x"cb" => c <= x"44";
				WHEN x"cc" => c <= x"75";
				WHEN x"cd" => c <= x"7e";
				WHEN x"ce" => c <= x"63";
				WHEN x"cf" => c <= x"68";  
				WHEN x"d0" => c <= x"b1";
				WHEN x"d1" => c <= x"ba";
				WHEN x"d2" => c <= x"a7";
				WHEN x"d3" => c <= x"ac";
				WHEN x"d4" => c <= x"9d";
				WHEN x"d5" => c <= x"96";
				WHEN x"d6" => c <= x"8b";
				WHEN x"d7" => c <= x"80";
				WHEN x"d8" => c <= x"e9";
				WHEN x"d9" => c <= x"e2";
				WHEN x"da" => c <= x"ff";
				WHEN x"db" => c <= x"f4";
				WHEN x"dc" => c <= x"c5";
				WHEN x"dd" => c <= x"ce";
				WHEN x"de" => c <= x"d3";
				WHEN x"df" => c <= x"d8"; 
				WHEN x"e0" => c <= x"7a";
				WHEN x"e1" => c <= x"71";
				WHEN x"e2" => c <= x"6c";
				WHEN x"e3" => c <= x"67";
				WHEN x"e4" => c <= x"56";
				WHEN x"e5" => c <= x"5d";
				WHEN x"e6" => c <= x"40";
				WHEN x"e7" => c <= x"4b";
				WHEN x"e8" => c <= x"22";
				WHEN x"e9" => c <= x"29";
				WHEN x"ea" => c <= x"34";
				WHEN x"eb" => c <= x"3f";
				WHEN x"ec" => c <= x"0e";
				WHEN x"ed" => c <= x"05";
				WHEN x"ee" => c <= x"18";
				WHEN x"ef" => c <= x"13";  
				WHEN x"f0" => c <= x"ca";
				WHEN x"f1" => c <= x"c1";
				WHEN x"f2" => c <= x"dc";
				WHEN x"f3" => c <= x"d7";
				WHEN x"f4" => c <= x"e6";
				WHEN x"f5" => c <= x"ed";
				WHEN x"f6" => c <= x"f0";
				WHEN x"f7" => c <= x"fb";
				WHEN x"f8" => c <= x"92";
				WHEN x"f9" => c <= x"99";
				WHEN x"fa" => c <= x"84";
				WHEN x"fb" => c <= x"8f";
				WHEN x"fc" => c <= x"be";
				WHEN x"fd" => c <= x"b5";
				WHEN x"fe" => c <= x"a8";
				WHEN x"ff" => c <= x"a3";  
				WHEN others => null;  
			END CASE; 
		WHEN x"13" =>
			CASE b IS
				WHEN x"00" => c <= x"00"; 
				WHEN x"01" => c <= x"0d"; 
				WHEN x"02" => c <= x"1a"; 
				WHEN x"03" => c <= x"17"; 
				WHEN x"04" => c <= x"34"; 
				WHEN x"05" => c <= x"39"; 
				WHEN x"06" => c <= x"2e"; 
				WHEN x"07" => c <= x"23"; 
				WHEN x"08" => c <= x"68"; 
				WHEN x"09" => c <= x"65"; 
				WHEN x"0a" => c <= x"72"; 
				WHEN x"0b" => c <= x"7f"; 
				WHEN x"0c" => c <= x"5c"; 
				WHEN x"0d" => c <= x"51"; 
				WHEN x"0e" => c <= x"46"; 
				WHEN x"0f" => c <= x"4b";  
				WHEN x"10" => c <= x"d0"; 
				WHEN x"11" => c <= x"dd"; 
				WHEN x"12" => c <= x"ca"; 
				WHEN x"13" => c <= x"c7"; 
				WHEN x"14" => c <= x"e4"; 
				WHEN x"15" => c <= x"e9"; 
				WHEN x"16" => c <= x"fe"; 
				WHEN x"17" => c <= x"f3"; 
				WHEN x"18" => c <= x"b8"; 
				WHEN x"19" => c <= x"b5"; 
				WHEN x"1a" => c <= x"a2"; 
				WHEN x"1b" => c <= x"af"; 
				WHEN x"1c" => c <= x"8c"; 
				WHEN x"1d" => c <= x"81"; 
				WHEN x"1e" => c <= x"96"; 
				WHEN x"1f" => c <= x"9b";
				WHEN x"20" => c <= x"bb";
				WHEN x"21" => c <= x"b6"; 
				WHEN x"22" => c <= x"a1"; 
				WHEN x"23" => c <= x"ac"; 
				WHEN x"24" => c <= x"8f"; 
				WHEN x"25" => c <= x"82"; 
				WHEN x"26" => c <= x"95"; 
				WHEN x"27" => c <= x"98"; 
				WHEN x"28" => c <= x"d3"; 
				WHEN x"29" => c <= x"de"; 
				WHEN x"2a" => c <= x"c9"; 
				WHEN x"2b" => c <= x"c4"; 
				WHEN x"2c" => c <= x"e7"; 
				WHEN x"2d" => c <= x"ea"; 
				WHEN x"2e" => c <= x"fd"; 
				WHEN x"2f" => c <= x"f0";  
				WHEN x"30" => c <= x"6b"; 
				WHEN x"31" => c <= x"66"; 
				WHEN x"32" => c <= x"71"; 
				WHEN x"33" => c <= x"7c"; 
				WHEN x"34" => c <= x"5f"; 
				WHEN x"35" => c <= x"52"; 
				WHEN x"36" => c <= x"45"; 
				WHEN x"37" => c <= x"48"; 
				WHEN x"38" => c <= x"03"; 
				WHEN x"39" => c <= x"0e"; 
				WHEN x"3a" => c <= x"19"; 
				WHEN x"3b" => c <= x"14"; 
				WHEN x"3c" => c <= x"37"; 
				WHEN x"3d" => c <= x"3a"; 
				WHEN x"3e" => c <= x"2d"; 
				WHEN x"3f" => c <= x"20";
				WHEN x"40" => c <= x"6d"; 
				WHEN x"41" => c <= x"60"; 
				WHEN x"42" => c <= x"77"; 
				WHEN x"43" => c <= x"7a"; 
				WHEN x"44" => c <= x"59"; 
				WHEN x"45" => c <= x"54"; 
				WHEN x"46" => c <= x"43"; 
				WHEN x"47" => c <= x"4e"; 
				WHEN x"48" => c <= x"05"; 
				WHEN x"49" => c <= x"08"; 
				WHEN x"4a" => c <= x"1f"; 
				WHEN x"4b" => c <= x"12"; 
				WHEN x"4c" => c <= x"31"; 
				WHEN x"4d" => c <= x"3c"; 
				WHEN x"4e" => c <= x"2b"; 
				WHEN x"4f" => c <= x"26";  
				WHEN x"50" => c <= x"bd";
				WHEN x"51" => c <= x"b0";
				WHEN x"52" => c <= x"a7";
				WHEN x"53" => c <= x"aa";
				WHEN x"54" => c <= x"89";
				WHEN x"55" => c <= x"84";
				WHEN x"56" => c <= x"93";
				WHEN x"57" => c <= x"9e";
				WHEN x"58" => c <= x"d5";
				WHEN x"59" => c <= x"d8";
				WHEN x"5a" => c <= x"cf";
				WHEN x"5b" => c <= x"c2";
				WHEN x"5c" => c <= x"e1";
				WHEN x"5d" => c <= x"ec";
				WHEN x"5e" => c <= x"fb";
				WHEN x"5f" => c <= x"f6"; 
				WHEN x"60" => c <= x"d6";
				WHEN x"61" => c <= x"db";
				WHEN x"62" => c <= x"cc";
				WHEN x"63" => c <= x"c1";
				WHEN x"64" => c <= x"e2";
				WHEN x"65" => c <= x"ef";
				WHEN x"66" => c <= x"f8";
				WHEN x"67" => c <= x"f5";
				WHEN x"68" => c <= x"be";
				WHEN x"69" => c <= x"b3";
				WHEN x"6a" => c <= x"a4";
				WHEN x"6b" => c <= x"a9";
				WHEN x"6c" => c <= x"8a";
				WHEN x"6d" => c <= x"87";
				WHEN x"6e" => c <= x"90";
				WHEN x"6f" => c <= x"9d";  
				WHEN x"70" => c <= x"06";
				WHEN x"71" => c <= x"0b";
				WHEN x"72" => c <= x"1c";
				WHEN x"73" => c <= x"11";
				WHEN x"74" => c <= x"32";
				WHEN x"75" => c <= x"3f";
				WHEN x"76" => c <= x"28";
				WHEN x"77" => c <= x"25";
				WHEN x"78" => c <= x"6e";
				WHEN x"79" => c <= x"63";
				WHEN x"7a" => c <= x"74";
				WHEN x"7b" => c <= x"79";
				WHEN x"7c" => c <= x"5a";
				WHEN x"7d" => c <= x"57";
				WHEN x"7e" => c <= x"40";
				WHEN x"7f" => c <= x"4d"; 
				WHEN x"80" => c <= x"da";
				WHEN x"81" => c <= x"d7";
				WHEN x"82" => c <= x"c0";
				WHEN x"83" => c <= x"cd";
				WHEN x"84" => c <= x"ee";
				WHEN x"85" => c <= x"e3";
				WHEN x"86" => c <= x"f4";
				WHEN x"87" => c <= x"f9";
				WHEN x"88" => c <= x"b2";
				WHEN x"89" => c <= x"bf";
				WHEN x"8a" => c <= x"a8";
				WHEN x"8b" => c <= x"a5";
				WHEN x"8c" => c <= x"86";
				WHEN x"8d" => c <= x"8b";
				WHEN x"8e" => c <= x"9c";
				WHEN x"8f" => c <= x"91";  
				WHEN x"90" => c <= x"0a";
				WHEN x"91" => c <= x"07";
				WHEN x"92" => c <= x"10";
				WHEN x"93" => c <= x"1d";
				WHEN x"94" => c <= x"3e";
				WHEN x"95" => c <= x"33";
				WHEN x"96" => c <= x"24";
				WHEN x"97" => c <= x"29";
				WHEN x"98" => c <= x"62";
				WHEN x"99" => c <= x"6f";
				WHEN x"9a" => c <= x"78";
				WHEN x"9b" => c <= x"75";
				WHEN x"9c" => c <= x"56";
				WHEN x"9d" => c <= x"5b";
				WHEN x"9e" => c <= x"4c";
				WHEN x"9f" => c <= x"41"; 
				WHEN x"a0" => c <= x"61";
				WHEN x"a1" => c <= x"6c";
				WHEN x"a2" => c <= x"7b";
				WHEN x"a3" => c <= x"76";
				WHEN x"a4" => c <= x"55";
				WHEN x"a5" => c <= x"58";
				WHEN x"a6" => c <= x"4f";
				WHEN x"a7" => c <= x"42";
				WHEN x"a8" => c <= x"09";
				WHEN x"a9" => c <= x"04";
				WHEN x"aa" => c <= x"13";
				WHEN x"ab" => c <= x"1e";
				WHEN x"ac" => c <= x"3d";
				WHEN x"ad" => c <= x"30";
				WHEN x"ae" => c <= x"27";
				WHEN x"af" => c <= x"2a";  
				WHEN x"b0" => c <= x"b1";
				WHEN x"b1" => c <= x"bc";
				WHEN x"b2" => c <= x"ab";
				WHEN x"b3" => c <= x"a6";
				WHEN x"b4" => c <= x"85";
				WHEN x"b5" => c <= x"88";
				WHEN x"b6" => c <= x"9f";
				WHEN x"b7" => c <= x"92";
				WHEN x"b8" => c <= x"d9";
				WHEN x"b9" => c <= x"d4";
				WHEN x"ba" => c <= x"c3";
				WHEN x"bb" => c <= x"ce";
				WHEN x"bc" => c <= x"ed";
				WHEN x"bd" => c <= x"e0";
				WHEN x"be" => c <= x"f7";
				WHEN x"bf" => c <= x"fa";
				WHEN x"c0" => c <= x"b7";
				WHEN x"c1" => c <= x"ba";
				WHEN x"c2" => c <= x"ad";
				WHEN x"c3" => c <= x"a0";
				WHEN x"c4" => c <= x"83";
				WHEN x"c5" => c <= x"8e";
				WHEN x"c6" => c <= x"99";
				WHEN x"c7" => c <= x"94";
				WHEN x"c8" => c <= x"df";
				WHEN x"c9" => c <= x"d2";
				WHEN x"ca" => c <= x"c5";
				WHEN x"cb" => c <= x"c8";
				WHEN x"cc" => c <= x"eb";
				WHEN x"cd" => c <= x"e6";
				WHEN x"ce" => c <= x"f1";
				WHEN x"cf" => c <= x"fc";  
				WHEN x"d0" => c <= x"67";
				WHEN x"d1" => c <= x"6a";
				WHEN x"d2" => c <= x"7d";
				WHEN x"d3" => c <= x"70";
				WHEN x"d4" => c <= x"53";
				WHEN x"d5" => c <= x"5e";
				WHEN x"d6" => c <= x"49";
				WHEN x"d7" => c <= x"44";
				WHEN x"d8" => c <= x"0f";
				WHEN x"d9" => c <= x"02";
				WHEN x"da" => c <= x"15";
				WHEN x"db" => c <= x"18";
				WHEN x"dc" => c <= x"3b";
				WHEN x"dd" => c <= x"36";
				WHEN x"de" => c <= x"21";
				WHEN x"df" => c <= x"2c"; 
				WHEN x"e0" => c <= x"0c";
				WHEN x"e1" => c <= x"01";
				WHEN x"e2" => c <= x"16";
				WHEN x"e3" => c <= x"1b";
				WHEN x"e4" => c <= x"38";
				WHEN x"e5" => c <= x"35";
				WHEN x"e6" => c <= x"22";
				WHEN x"e7" => c <= x"2f";
				WHEN x"e8" => c <= x"64";
				WHEN x"e9" => c <= x"69";
				WHEN x"ea" => c <= x"7e";
				WHEN x"eb" => c <= x"73";
				WHEN x"ec" => c <= x"50";
				WHEN x"ed" => c <= x"5d";
				WHEN x"ee" => c <= x"4a";
				WHEN x"ef" => c <= x"47";  
				WHEN x"f0" => c <= x"dc";
				WHEN x"f1" => c <= x"d1";
				WHEN x"f2" => c <= x"c6";
				WHEN x"f3" => c <= x"cb";
				WHEN x"f4" => c <= x"e8";
				WHEN x"f5" => c <= x"e5";
				WHEN x"f6" => c <= x"f2";
				WHEN x"f7" => c <= x"ff";
				WHEN x"f8" => c <= x"b4";
				WHEN x"f9" => c <= x"b9";
				WHEN x"fa" => c <= x"ae";
				WHEN x"fb" => c <= x"a3";
				WHEN x"fc" => c <= x"80";
				WHEN x"fd" => c <= x"8d";
				WHEN x"fe" => c <= x"9a";
				WHEN x"ff" => c <= x"97";  
				WHEN others => null;  
			END CASE; 
		WHEN x"14" =>
			CASE b IS
				WHEN x"00" => c <= x"00"; 
				WHEN x"01" => c <= x"0e"; 
				WHEN x"02" => c <= x"1c"; 
				WHEN x"03" => c <= x"12"; 
				WHEN x"04" => c <= x"38"; 
				WHEN x"05" => c <= x"36"; 
				WHEN x"06" => c <= x"24"; 
				WHEN x"07" => c <= x"2a"; 
				WHEN x"08" => c <= x"70"; 
				WHEN x"09" => c <= x"7e"; 
				WHEN x"0a" => c <= x"6c"; 
				WHEN x"0b" => c <= x"62"; 
				WHEN x"0c" => c <= x"48"; 
				WHEN x"0d" => c <= x"46"; 
				WHEN x"0e" => c <= x"54"; 
				WHEN x"0f" => c <= x"5a";  
				WHEN x"10" => c <= x"e0"; 
				WHEN x"11" => c <= x"ee"; 
				WHEN x"12" => c <= x"fc"; 
				WHEN x"13" => c <= x"f2"; 
				WHEN x"14" => c <= x"d8"; 
				WHEN x"15" => c <= x"d6"; 
				WHEN x"16" => c <= x"c4"; 
				WHEN x"17" => c <= x"ca"; 
				WHEN x"18" => c <= x"90"; 
				WHEN x"19" => c <= x"9e"; 
				WHEN x"1a" => c <= x"8c"; 
				WHEN x"1b" => c <= x"82"; 
				WHEN x"1c" => c <= x"a8"; 
				WHEN x"1d" => c <= x"a6"; 
				WHEN x"1e" => c <= x"b4"; 
				WHEN x"1f" => c <= x"ba";
				WHEN x"20" => c <= x"db";
				WHEN x"21" => c <= x"d5"; 
				WHEN x"22" => c <= x"c7"; 
				WHEN x"23" => c <= x"c9"; 
				WHEN x"24" => c <= x"e3"; 
				WHEN x"25" => c <= x"ed"; 
				WHEN x"26" => c <= x"ff"; 
				WHEN x"27" => c <= x"f1"; 
				WHEN x"28" => c <= x"ab"; 
				WHEN x"29" => c <= x"a5"; 
				WHEN x"2a" => c <= x"b7"; 
				WHEN x"2b" => c <= x"b9"; 
				WHEN x"2c" => c <= x"93"; 
				WHEN x"2d" => c <= x"9d"; 
				WHEN x"2e" => c <= x"8f"; 
				WHEN x"2f" => c <= x"81";  
				WHEN x"30" => c <= x"3b"; 
				WHEN x"31" => c <= x"35"; 
				WHEN x"32" => c <= x"27"; 
				WHEN x"33" => c <= x"29"; 
				WHEN x"34" => c <= x"03"; 
				WHEN x"35" => c <= x"0d"; 
				WHEN x"36" => c <= x"1f"; 
				WHEN x"37" => c <= x"11"; 
				WHEN x"38" => c <= x"4b"; 
				WHEN x"39" => c <= x"45"; 
				WHEN x"3a" => c <= x"57"; 
				WHEN x"3b" => c <= x"59"; 
				WHEN x"3c" => c <= x"73"; 
				WHEN x"3d" => c <= x"7d"; 
				WHEN x"3e" => c <= x"6f"; 
				WHEN x"3f" => c <= x"61";
				WHEN x"40" => c <= x"ad"; 
				WHEN x"41" => c <= x"a3"; 
				WHEN x"42" => c <= x"b1"; 
				WHEN x"43" => c <= x"bf"; 
				WHEN x"44" => c <= x"95"; 
				WHEN x"45" => c <= x"9b"; 
				WHEN x"46" => c <= x"89"; 
				WHEN x"47" => c <= x"87"; 
				WHEN x"48" => c <= x"dd"; 
				WHEN x"49" => c <= x"d3"; 
				WHEN x"4a" => c <= x"c1"; 
				WHEN x"4b" => c <= x"cf"; 
				WHEN x"4c" => c <= x"e5"; 
				WHEN x"4d" => c <= x"eb"; 
				WHEN x"4e" => c <= x"f9"; 
				WHEN x"4f" => c <= x"f7";  
				WHEN x"50" => c <= x"4d";
				WHEN x"51" => c <= x"43";
				WHEN x"52" => c <= x"51";
				WHEN x"53" => c <= x"5f";
				WHEN x"54" => c <= x"75";
				WHEN x"55" => c <= x"7b";
				WHEN x"56" => c <= x"69";
				WHEN x"57" => c <= x"67";
				WHEN x"58" => c <= x"3d";
				WHEN x"59" => c <= x"33";
				WHEN x"5a" => c <= x"21";
				WHEN x"5b" => c <= x"2f";
				WHEN x"5c" => c <= x"05";
				WHEN x"5d" => c <= x"0b";
				WHEN x"5e" => c <= x"19";
				WHEN x"5f" => c <= x"17"; 
				WHEN x"60" => c <= x"76";
				WHEN x"61" => c <= x"78";
				WHEN x"62" => c <= x"6a";
				WHEN x"63" => c <= x"64";
				WHEN x"64" => c <= x"4e";
				WHEN x"65" => c <= x"40";
				WHEN x"66" => c <= x"52";
				WHEN x"67" => c <= x"5c";
				WHEN x"68" => c <= x"06";
				WHEN x"69" => c <= x"08";
				WHEN x"6a" => c <= x"1a";
				WHEN x"6b" => c <= x"14";
				WHEN x"6c" => c <= x"3e";
				WHEN x"6d" => c <= x"30";
				WHEN x"6e" => c <= x"22";
				WHEN x"6f" => c <= x"2c";  
				WHEN x"70" => c <= x"96";
				WHEN x"71" => c <= x"98";
				WHEN x"72" => c <= x"8a";
				WHEN x"73" => c <= x"84";
				WHEN x"74" => c <= x"ae";
				WHEN x"75" => c <= x"a0";
				WHEN x"76" => c <= x"b2";
				WHEN x"77" => c <= x"bc";
				WHEN x"78" => c <= x"e6";
				WHEN x"79" => c <= x"e8";
				WHEN x"7a" => c <= x"fa";
				WHEN x"7b" => c <= x"f4";
				WHEN x"7c" => c <= x"de";
				WHEN x"7d" => c <= x"d0";
				WHEN x"7e" => c <= x"c2";
				WHEN x"7f" => c <= x"cc"; 
				WHEN x"80" => c <= x"41";
				WHEN x"81" => c <= x"4f";
				WHEN x"82" => c <= x"5d";
				WHEN x"83" => c <= x"53";
				WHEN x"84" => c <= x"79";
				WHEN x"85" => c <= x"77";
				WHEN x"86" => c <= x"65";
				WHEN x"87" => c <= x"6b";
				WHEN x"88" => c <= x"31";
				WHEN x"89" => c <= x"3f";
				WHEN x"8a" => c <= x"2d";
				WHEN x"8b" => c <= x"23";
				WHEN x"8c" => c <= x"09";
				WHEN x"8d" => c <= x"07";
				WHEN x"8e" => c <= x"15";
				WHEN x"8f" => c <= x"1b";  
				WHEN x"90" => c <= x"a1";
				WHEN x"91" => c <= x"af";
				WHEN x"92" => c <= x"bd";
				WHEN x"93" => c <= x"b3";
				WHEN x"94" => c <= x"99";
				WHEN x"95" => c <= x"97";
				WHEN x"96" => c <= x"85";
				WHEN x"97" => c <= x"8b";
				WHEN x"98" => c <= x"d1";
				WHEN x"99" => c <= x"df";
				WHEN x"9a" => c <= x"cd";
				WHEN x"9b" => c <= x"c3";
				WHEN x"9c" => c <= x"e9";
				WHEN x"9d" => c <= x"e7";
				WHEN x"9e" => c <= x"f5";
				WHEN x"9f" => c <= x"fb"; 
				WHEN x"a0" => c <= x"9a";
				WHEN x"a1" => c <= x"94";
				WHEN x"a2" => c <= x"86";
				WHEN x"a3" => c <= x"88";
				WHEN x"a4" => c <= x"a2";
				WHEN x"a5" => c <= x"ac";
				WHEN x"a6" => c <= x"be";
				WHEN x"a7" => c <= x"b0";
				WHEN x"a8" => c <= x"ea";
				WHEN x"a9" => c <= x"e4";
				WHEN x"aa" => c <= x"f6";
				WHEN x"ab" => c <= x"f8";
				WHEN x"ac" => c <= x"d2";
				WHEN x"ad" => c <= x"dc";
				WHEN x"ae" => c <= x"ce";
				WHEN x"af" => c <= x"c0";  
				WHEN x"b0" => c <= x"7a";
				WHEN x"b1" => c <= x"74";
				WHEN x"b2" => c <= x"66";
				WHEN x"b3" => c <= x"68";
				WHEN x"b4" => c <= x"42";
				WHEN x"b5" => c <= x"4c";
				WHEN x"b6" => c <= x"5e";
				WHEN x"b7" => c <= x"50";
				WHEN x"b8" => c <= x"0a";
				WHEN x"b9" => c <= x"04";
				WHEN x"ba" => c <= x"16";
				WHEN x"bb" => c <= x"18";
				WHEN x"bc" => c <= x"32";
				WHEN x"bd" => c <= x"3c";
				WHEN x"be" => c <= x"2e";
				WHEN x"bf" => c <= x"20";
				WHEN x"c0" => c <= x"ec";
				WHEN x"c1" => c <= x"e2";
				WHEN x"c2" => c <= x"f0";
				WHEN x"c3" => c <= x"fe";
				WHEN x"c4" => c <= x"d4";
				WHEN x"c5" => c <= x"da";
				WHEN x"c6" => c <= x"c8";
				WHEN x"c7" => c <= x"c6";
				WHEN x"c8" => c <= x"9c";
				WHEN x"c9" => c <= x"92";
				WHEN x"ca" => c <= x"80";
				WHEN x"cb" => c <= x"8e";
				WHEN x"cc" => c <= x"a4";
				WHEN x"cd" => c <= x"aa";
				WHEN x"ce" => c <= x"b8";
				WHEN x"cf" => c <= x"b6";  
				WHEN x"d0" => c <= x"0c";
				WHEN x"d1" => c <= x"02";
				WHEN x"d2" => c <= x"10";
				WHEN x"d3" => c <= x"1e";
				WHEN x"d4" => c <= x"34";
				WHEN x"d5" => c <= x"3a";
				WHEN x"d6" => c <= x"28";
				WHEN x"d7" => c <= x"26";
				WHEN x"d8" => c <= x"7c";
				WHEN x"d9" => c <= x"72";
				WHEN x"da" => c <= x"60";
				WHEN x"db" => c <= x"6e";
				WHEN x"dc" => c <= x"44";
				WHEN x"dd" => c <= x"4a";
				WHEN x"de" => c <= x"58";
				WHEN x"df" => c <= x"56"; 
				WHEN x"e0" => c <= x"37";
				WHEN x"e1" => c <= x"39";
				WHEN x"e2" => c <= x"2b";
				WHEN x"e3" => c <= x"25";
				WHEN x"e4" => c <= x"0f";
				WHEN x"e5" => c <= x"01";
				WHEN x"e6" => c <= x"13";
				WHEN x"e7" => c <= x"1d";
				WHEN x"e8" => c <= x"47";
				WHEN x"e9" => c <= x"49";
				WHEN x"ea" => c <= x"5b";
				WHEN x"eb" => c <= x"55";
				WHEN x"ec" => c <= x"7f";
				WHEN x"ed" => c <= x"71";
				WHEN x"ee" => c <= x"63";
				WHEN x"ef" => c <= x"6d";  
				WHEN x"f0" => c <= x"d7";
				WHEN x"f1" => c <= x"d9";
				WHEN x"f2" => c <= x"cb";
				WHEN x"f3" => c <= x"c5";
				WHEN x"f4" => c <= x"ef";
				WHEN x"f5" => c <= x"e1";
				WHEN x"f6" => c <= x"f3";
				WHEN x"f7" => c <= x"fd";
				WHEN x"f8" => c <= x"a7";
				WHEN x"f9" => c <= x"a9";
				WHEN x"fa" => c <= x"bb";
				WHEN x"fb" => c <= x"b5";
				WHEN x"fc" => c <= x"9f";
				WHEN x"fd" => c <= x"91";
				WHEN x"fe" => c <= x"83";
				WHEN x"ff" => c <= x"8d";  
				WHEN others => null;  
			END CASE; 
			
			WHEN others => null; 
		END CASE;
  END PROCESS find;
END rtl;

