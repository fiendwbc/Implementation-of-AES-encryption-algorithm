LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_ARITH.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE work.ALL;
USE work.type_pkg.ALL;

ENTITY sbox_lookup IS
  PORT(a: IN SLV_8; b: OUT SLV_8);
END sbox_lookup;
ARCHITECTURE rtl OF sbox_lookup IS
BEGIN
   P0: PROCESS(a)
	BEGIN 
	CASE a IS   
		WHEN x"00" => b <= x"63"; 
		WHEN x"01" => b <= x"7c"; 
		WHEN x"02" => b <= x"77"; 
		WHEN x"03" => b <= x"7b"; 
		WHEN x"04" => b <= x"f2"; 
		WHEN x"05" => b <= x"6b"; 
		WHEN x"06" => b <= x"6f"; 
		WHEN x"07" => b <= x"c5"; 
		WHEN x"08" => b <= x"30"; 
		WHEN x"09" => b <= x"01"; 
		WHEN x"0a" => b <= x"67"; 
		WHEN x"0b" => b <= x"2b"; 
		WHEN x"0c" => b <= x"fe"; 
		WHEN x"0d" => b <= x"d7"; 
		WHEN x"0e" => b <= x"ab"; 
		WHEN x"0f" => b <= x"76";  
		WHEN x"10" => b <= x"ca"; 
		WHEN x"11" => b <= x"82"; 
		WHEN x"12" => b <= x"c9"; 
		WHEN x"13" => b <= x"7d"; 
		WHEN x"14" => b <= x"fa"; 
		WHEN x"15" => b <= x"59"; 
		WHEN x"16" => b <= x"47"; 
		WHEN x"17" => b <= x"f0"; 
		WHEN x"18" => b <= x"ad"; 
		WHEN x"19" => b <= x"d4"; 
		WHEN x"1a" => b <= x"a2"; 
		WHEN x"1b" => b <= x"af"; 
		WHEN x"1c" => b <= x"9c"; 
		WHEN x"1d" => b <= x"a4"; 
		WHEN x"1e" => b <= x"72"; 
		WHEN x"1f" => b <= x"c0";
		WHEN x"20" => b <= x"b7";
		WHEN x"21" => b <= x"fd"; 
		WHEN x"22" => b <= x"93"; 
		WHEN x"23" => b <= x"26"; 
		WHEN x"24" => b <= x"36"; 
		WHEN x"25" => b <= x"3f"; 
		WHEN x"26" => b <= x"f7"; 
		WHEN x"27" => b <= x"cc"; 
		WHEN x"28" => b <= x"34"; 
		WHEN x"29" => b <= x"a5"; 
		WHEN x"2a" => b <= x"e5"; 
		WHEN x"2b" => b <= x"f1"; 
		WHEN x"2c" => b <= x"71"; 
		WHEN x"2d" => b <= x"d8"; 
		WHEN x"2e" => b <= x"31"; 
		WHEN x"2f" => b <= x"15";  
		WHEN x"30" => b <= x"04"; 
		WHEN x"31" => b <= x"c7"; 
				WHEN x"32" => b <= x"23"; 
				WHEN x"33" => b <= x"c3"; 
				WHEN x"34" => b <= x"18"; 
				WHEN x"35" => b <= x"96"; 
				WHEN x"36" => b <= x"05"; 
				WHEN x"37" => b <= x"9a"; 
				WHEN x"38" => b <= x"07"; 
				WHEN x"39" => b <= x"12"; 
				WHEN x"3a" => b <= x"80"; 
				WHEN x"3b" => b <= x"e2"; 
				WHEN x"3c" => b <= x"eb"; 
				WHEN x"3d" => b <= x"27"; 
				WHEN x"3e" => b <= x"b2"; 
				WHEN x"3f" => b <= x"75";
				WHEN x"40" => b <= x"09"; 
				WHEN x"41" => b <= x"83"; 
				WHEN x"42" => b <= x"2c"; 
				WHEN x"43" => b <= x"1a"; 
				WHEN x"44" => b <= x"1b"; 
				WHEN x"45" => b <= x"6e"; 
				WHEN x"46" => b <= x"5a"; 
				WHEN x"47" => b <= x"a0"; 
				WHEN x"48" => b <= x"52"; 
				WHEN x"49" => b <= x"3b"; 
				WHEN x"4a" => b <= x"d6"; 
				WHEN x"4b" => b <= x"b3"; 
				WHEN x"4c" => b <= x"29"; 
				WHEN x"4d" => b <= x"e3"; 
				WHEN x"4e" => b <= x"2f"; 
				WHEN x"4f" => b <= x"84";  
				 
				WHEN x"50" => b <= x"53";
				WHEN x"51" => b <= x"d1";
				WHEN x"52" => b <= x"00";
				WHEN x"53" => b <= x"ed";
				WHEN x"54" => b <= x"20";
				WHEN x"55" => b <= x"fc";
				WHEN x"56" => b <= x"b1";
				WHEN x"57" => b <= x"5b";
				WHEN x"58" => b <= x"6a";
				WHEN x"59" => b <= x"cb";
				WHEN x"5a" => b <= x"be";
				WHEN x"5b" => b <= x"39";
				WHEN x"5c" => b <= x"4a";
				WHEN x"5d" => b <= x"4c";
				WHEN x"5e" => b <= x"58";
				WHEN x"5f" => b <= x"cf"; 
				WHEN x"60" => b <= x"d0";
				WHEN x"61" => b <= x"ef";
				WHEN x"62" => b <= x"aa";
				WHEN x"63" => b <= x"fb";
				WHEN x"64" => b <= x"43";
				WHEN x"65" => b <= x"4d";
				WHEN x"66" => b <= x"33";
				WHEN x"67" => b <= x"85";
				WHEN x"68" => b <= x"45";
				WHEN x"69" => b <= x"f9";
				WHEN x"6a" => b <= x"02";
				WHEN x"6b" => b <= x"7f";
				WHEN x"6c" => b <= x"50";
				WHEN x"6d" => b <= x"3c";
				WHEN x"6e" => b <= x"9f";
				WHEN x"6f" => b <= x"a8";  
				WHEN x"70" => b <= x"51";
				WHEN x"71" => b <= x"a3";
				WHEN x"72" => b <= x"40";
				WHEN x"73" => b <= x"8f";
				WHEN x"74" => b <= x"92";
				WHEN x"75" => b <= x"9d";
				WHEN x"76" => b <= x"38";
				WHEN x"77" => b <= x"f5";
				WHEN x"78" => b <= x"bc";
				WHEN x"79" => b <= x"b6";
				WHEN x"7a" => b <= x"da";
				WHEN x"7b" => b <= x"21";
				WHEN x"7c" => b <= x"10";
				WHEN x"7d" => b <= x"ff";
				WHEN x"7e" => b <= x"f3";
				WHEN x"7f" => b <= x"d2"; 
				WHEN x"80" => b <= x"cd";
				WHEN x"81" => b <= x"0c";
				WHEN x"82" => b <= x"13";
				WHEN x"83" => b <= x"ec";
				WHEN x"84" => b <= x"5f";
				WHEN x"85" => b <= x"97";
				WHEN x"86" => b <= x"44";
				WHEN x"87" => b <= x"17";
				WHEN x"88" => b <= x"c4";
				WHEN x"89" => b <= x"a7";
				WHEN x"8a" => b <= x"7e";
				WHEN x"8b" => b <= x"3d";
				WHEN x"8c" => b <= x"64";
				WHEN x"8d" => b <= x"5d";
				WHEN x"8e" => b <= x"19";
				WHEN x"8f" => b <= x"73";  
				WHEN x"90" => b <= x"60";
				WHEN x"91" => b <= x"81";
				WHEN x"92" => b <= x"4f";
				WHEN x"93" => b <= x"dc";
				WHEN x"94" => b <= x"22";
				WHEN x"95" => b <= x"2a";
				WHEN x"96" => b <= x"90";
				WHEN x"97" => b <= x"88";
				WHEN x"98" => b <= x"46";
				WHEN x"99" => b <= x"ee";
				WHEN x"9a" => b <= x"b8";
				WHEN x"9b" => b <= x"14";
				WHEN x"9c" => b <= x"de";
				WHEN x"9d" => b <= x"5e";
				WHEN x"9e" => b <= x"0b";
				WHEN x"9f" => b <= x"db"; 
				WHEN x"a0" => b <= x"e0";
				WHEN x"a1" => b <= x"32";
				WHEN x"a2" => b <= x"3a";
				WHEN x"a3" => b <= x"0a";
				WHEN x"a4" => b <= x"49";
				WHEN x"a5" => b <= x"06";
				WHEN x"a6" => b <= x"24";
				WHEN x"a7" => b <= x"5c";
				WHEN x"a8" => b <= x"c2";
				WHEN x"a9" => b <= x"d3";
				WHEN x"aa" => b <= x"ac";
				WHEN x"ab" => b <= x"62";
				WHEN x"ac" => b <= x"91";
				WHEN x"ad" => b <= x"95";
				WHEN x"ae" => b <= x"e4";
				WHEN x"af" => b <= x"79";  
				WHEN x"b0" => b <= x"e7";
				WHEN x"b1" => b <= x"c8";
				WHEN x"b2" => b <= x"37";
				WHEN x"b3" => b <= x"6d";
				WHEN x"b4" => b <= x"8d";
				WHEN x"b5" => b <= x"d5";
				WHEN x"b6" => b <= x"4e";
				WHEN x"b7" => b <= x"a9";
				WHEN x"b8" => b <= x"6c";
				WHEN x"b9" => b <= x"56";
				WHEN x"ba" => b <= x"f4";
				WHEN x"bb" => b <= x"ea";
				WHEN x"bc" => b <= x"65";
				WHEN x"bd" => b <= x"7a";
				WHEN x"be" => b <= x"ae";
				WHEN x"bf" => b <= x"08";
				WHEN x"c0" => b <= x"ba";
				WHEN x"c1" => b <= x"78";
				WHEN x"c2" => b <= x"25";
				WHEN x"c3" => b <= x"2e";
				WHEN x"c4" => b <= x"1c";
				WHEN x"c5" => b <= x"a6";
				WHEN x"c6" => b <= x"b4";
				WHEN x"c7" => b <= x"c6";
				WHEN x"c8" => b <= x"e8";
				WHEN x"c9" => b <= x"dd";
				WHEN x"ca" => b <= x"74";
				WHEN x"cb" => b <= x"1f";
				WHEN x"cc" => b <= x"4b";
				WHEN x"cd" => b <= x"bd";
				WHEN x"ce" => b <= x"8b";
				WHEN x"cf" => b <= x"8a";  
				WHEN x"d0" => b <= x"70";
				WHEN x"d1" => b <= x"3e";
				WHEN x"d2" => b <= x"b5";
				WHEN x"d3" => b <= x"66";
				WHEN x"d4" => b <= x"48";
				WHEN x"d5" => b <= x"03";
				WHEN x"d6" => b <= x"f6";
				WHEN x"d7" => b <= x"0e";
				WHEN x"d8" => b <= x"61";
				WHEN x"d9" => b <= x"35";
				WHEN x"da" => b <= x"57";
				WHEN x"db" => b <= x"b9";
				WHEN x"dc" => b <= x"86";
				WHEN x"dd" => b <= x"c1";
				WHEN x"de" => b <= x"1d";
				WHEN x"df" => b <= x"9e"; 
				WHEN x"e0" => b <= x"e1";
				WHEN x"e1" => b <= x"f8";
				WHEN x"e2" => b <= x"98";
				WHEN x"e3" => b <= x"11";
				WHEN x"e4" => b <= x"69";
				WHEN x"e5" => b <= x"d9";
				WHEN x"e6" => b <= x"8e";
				WHEN x"e7" => b <= x"94";
				WHEN x"e8" => b <= x"9b";
				WHEN x"e9" => b <= x"1e";
				WHEN x"ea" => b <= x"87";
				WHEN x"eb" => b <= x"e9";
				WHEN x"ec" => b <= x"ce";
				WHEN x"ed" => b <= x"55";
				WHEN x"ee" => b <= x"28";
				WHEN x"ef" => b <= x"df";  
				WHEN x"f0" => b <= x"8c";
				WHEN x"f1" => b <= x"a1";
				WHEN x"f2" => b <= x"89";
				WHEN x"f3" => b <= x"0d";
				WHEN x"f4" => b <= x"bf";
				WHEN x"f5" => b <= x"e6";
				WHEN x"f6" => b <= x"42";
				WHEN x"f7" => b <= x"68";
				WHEN x"f8" => b <= x"41";
				WHEN x"f9" => b <= x"99";
				WHEN x"fa" => b <= x"2d";
				WHEN x"fb" => b <= x"0f";
				WHEN x"fc" => b <= x"b0";
				WHEN x"fd" => b <= x"54";
				WHEN x"fe" => b <= x"bb";
				WHEN x"ff" => b <= x"16";  
				WHEN others => null;  
			END CASE;   
		END PROCESS P0;
END rtl;




