LIBRARY IEEE; 
USE IEEE.STD_LOGIC_1164.ALL; 
USE work.ALL;
USE work.type_pkg.ALL;

ENTITY states_substitute_process IS
  PORT(state: IN STATE_ARRAY; 
  num: IN INTEGER;
  state_after_sub: OUT STATE_ARRAY);
END states_substitute_process;
  
ARCHITECTURE rtl OF states_substitute_process IS
  COMPONENT sbox_lookup
      PORT(a: IN SLV_8; b: OUT SLV_8);
  END COMPONENT;
 -- SIGNAL cWord: SLV_8;
 -- SIGNAL b: SLV_8;
 -- SIGNAL cIndex: INTEGER :=0;
 -- SIGNAL t: STATE_ARRAY;
BEGIN
  find:PROCESS(num)
    BEGIN
      FOR I IN 0 TO 15 LOOP
--        sbox_lookup PORT MAP(state(I), t(I));
	     	CASE state(I) IS   
			WHEN x"00" => state_after_sub(I) <= x"63"; 
			WHEN x"01" => state_after_sub(I) <= x"7c"; 
			WHEN x"02" => state_after_sub(I) <= x"77"; 
			WHEN x"03" => state_after_sub(I) <= x"7b"; 
			WHEN x"04" => state_after_sub(I) <= x"f2"; 
			WHEN x"05" => state_after_sub(I) <= x"6b"; 
			WHEN x"06" => state_after_sub(I) <= x"6f"; 
			WHEN x"07" => state_after_sub(I) <= x"c5"; 
			WHEN x"08" => state_after_sub(I) <= x"30"; 
			WHEN x"09" => state_after_sub(I) <= x"01"; 
			WHEN x"0a" => state_after_sub(I) <= x"67"; 
			WHEN x"0b" => state_after_sub(I) <= x"2b"; 
			WHEN x"0c" => state_after_sub(I) <= x"fe"; 
			WHEN x"0d" => state_after_sub(I) <= x"d7"; 
			WHEN x"0e" => state_after_sub(I) <= x"ab"; 
			WHEN x"0f" => state_after_sub(I) <= x"76";  
			WHEN x"10" => state_after_sub(I) <= x"ca"; 
			WHEN x"11" => state_after_sub(I) <= x"82"; 
			WHEN x"12" => state_after_sub(I) <= x"c9"; 
			WHEN x"13" => state_after_sub(I) <= x"7d"; 
			WHEN x"14" => state_after_sub(I) <= x"fa"; 
			WHEN x"15" => state_after_sub(I) <= x"59"; 
			WHEN x"16" => state_after_sub(I) <= x"47"; 
			WHEN x"17" => state_after_sub(I) <= x"f0"; 
			WHEN x"18" => state_after_sub(I) <= x"ad"; 
			WHEN x"19" => state_after_sub(I) <= x"d4"; 
			WHEN x"1a" => state_after_sub(I) <= x"a2"; 
			WHEN x"1b" => state_after_sub(I) <= x"af"; 
			WHEN x"1c" => state_after_sub(I) <= x"9c"; 
			WHEN x"1d" => state_after_sub(I) <= x"a4"; 
			WHEN x"1e" => state_after_sub(I) <= x"72"; 
			WHEN x"1f" => state_after_sub(I) <= x"c0";
			WHEN x"20" => state_after_sub(I) <= x"b7";
			WHEN x"21" => state_after_sub(I) <= x"fd"; 
			WHEN x"22" => state_after_sub(I) <= x"93"; 
			WHEN x"23" => state_after_sub(I) <= x"26"; 
			WHEN x"24" => state_after_sub(I) <= x"36"; 
			WHEN x"25" => state_after_sub(I) <= x"3f"; 
			WHEN x"26" => state_after_sub(I) <= x"f7"; 
			WHEN x"27" => state_after_sub(I) <= x"cc"; 
			WHEN x"28" => state_after_sub(I) <= x"34"; 
			WHEN x"29" => state_after_sub(I) <= x"a5"; 
			WHEN x"2a" => state_after_sub(I) <= x"e5"; 
			WHEN x"2b" => state_after_sub(I) <= x"f1"; 
			WHEN x"2c" => state_after_sub(I) <= x"71"; 
			WHEN x"2d" => state_after_sub(I) <= x"d8"; 
			WHEN x"2e" => state_after_sub(I) <= x"31"; 
			WHEN x"2f" => state_after_sub(I) <= x"15";  
			WHEN x"30" => state_after_sub(I) <= x"04"; 
			WHEN x"31" => state_after_sub(I) <= x"c7"; 
					WHEN x"32" => state_after_sub(I) <= x"23"; 
					WHEN x"33" => state_after_sub(I) <= x"c3"; 
					WHEN x"34" => state_after_sub(I) <= x"18"; 
					WHEN x"35" => state_after_sub(I) <= x"96"; 
					WHEN x"36" => state_after_sub(I) <= x"05"; 
					WHEN x"37" => state_after_sub(I) <= x"9a"; 
					WHEN x"38" => state_after_sub(I) <= x"07"; 
					WHEN x"39" => state_after_sub(I) <= x"12"; 
					WHEN x"3a" => state_after_sub(I) <= x"80"; 
					WHEN x"3b" => state_after_sub(I) <= x"e2"; 
					WHEN x"3c" => state_after_sub(I) <= x"eb"; 
					WHEN x"3d" => state_after_sub(I) <= x"27"; 
					WHEN x"3e" => state_after_sub(I) <= x"b2"; 
					WHEN x"3f" => state_after_sub(I) <= x"75";
					WHEN x"40" => state_after_sub(I) <= x"09"; 
					WHEN x"41" => state_after_sub(I) <= x"83"; 
					WHEN x"42" => state_after_sub(I) <= x"2c"; 
					WHEN x"43" => state_after_sub(I) <= x"1a"; 
					WHEN x"44" => state_after_sub(I) <= x"1b"; 
					WHEN x"45" => state_after_sub(I) <= x"6e"; 
					WHEN x"46" => state_after_sub(I) <= x"5a"; 
					WHEN x"47" => state_after_sub(I) <= x"a0"; 
					WHEN x"48" => state_after_sub(I) <= x"52"; 
					WHEN x"49" => state_after_sub(I) <= x"3b"; 
					WHEN x"4a" => state_after_sub(I) <= x"d6"; 
					WHEN x"4b" => state_after_sub(I) <= x"b3"; 
					WHEN x"4c" => state_after_sub(I) <= x"29"; 
					WHEN x"4d" => state_after_sub(I) <= x"e3"; 
					WHEN x"4e" => state_after_sub(I) <= x"2f"; 
					WHEN x"4f" => state_after_sub(I) <= x"84";  
					 
					WHEN x"50" => state_after_sub(I) <= x"53";
					WHEN x"51" => state_after_sub(I) <= x"d1";
					WHEN x"52" => state_after_sub(I) <= x"00";
					WHEN x"53" => state_after_sub(I) <= x"ed";
					WHEN x"54" => state_after_sub(I) <= x"20";
					WHEN x"55" => state_after_sub(I) <= x"fc";
					WHEN x"56" => state_after_sub(I) <= x"b1";
					WHEN x"57" => state_after_sub(I) <= x"5b";
					WHEN x"58" => state_after_sub(I) <= x"6a";
					WHEN x"59" => state_after_sub(I) <= x"cb";
					WHEN x"5a" => state_after_sub(I) <= x"be";
					WHEN x"5b" => state_after_sub(I) <= x"39";
					WHEN x"5c" => state_after_sub(I) <= x"4a";
					WHEN x"5d" => state_after_sub(I) <= x"4c";
					WHEN x"5e" => state_after_sub(I) <= x"58";
					WHEN x"5f" => state_after_sub(I) <= x"cf"; 
					WHEN x"60" => state_after_sub(I) <= x"d0";
					WHEN x"61" => state_after_sub(I) <= x"ef";
					WHEN x"62" => state_after_sub(I) <= x"aa";
					WHEN x"63" => state_after_sub(I) <= x"fb";
					WHEN x"64" => state_after_sub(I) <= x"43";
					WHEN x"65" => state_after_sub(I) <= x"4d";
					WHEN x"66" => state_after_sub(I) <= x"33";
					WHEN x"67" => state_after_sub(I) <= x"85";
					WHEN x"68" => state_after_sub(I) <= x"45";
					WHEN x"69" => state_after_sub(I) <= x"f9";
					WHEN x"6a" => state_after_sub(I) <= x"02";
					WHEN x"6b" => state_after_sub(I) <= x"7f";
					WHEN x"6c" => state_after_sub(I) <= x"50";
					WHEN x"6d" => state_after_sub(I) <= x"3c";
					WHEN x"6e" => state_after_sub(I) <= x"9f";
					WHEN x"6f" => state_after_sub(I) <= x"a8";  
					WHEN x"70" => state_after_sub(I) <= x"51";
					WHEN x"71" => state_after_sub(I) <= x"a3";
					WHEN x"72" => state_after_sub(I) <= x"40";
					WHEN x"73" => state_after_sub(I) <= x"8f";
					WHEN x"74" => state_after_sub(I) <= x"92";
					WHEN x"75" => state_after_sub(I) <= x"9d";
					WHEN x"76" => state_after_sub(I) <= x"38";
					WHEN x"77" => state_after_sub(I) <= x"f5";
					WHEN x"78" => state_after_sub(I) <= x"bc";
					WHEN x"79" => state_after_sub(I) <= x"b6";
					WHEN x"7a" => state_after_sub(I) <= x"da";
					WHEN x"7b" => state_after_sub(I) <= x"21";
					WHEN x"7c" => state_after_sub(I) <= x"10";
					WHEN x"7d" => state_after_sub(I) <= x"ff";
					WHEN x"7e" => state_after_sub(I) <= x"f3";
					WHEN x"7f" => state_after_sub(I) <= x"d2"; 
					WHEN x"80" => state_after_sub(I) <= x"cd";
					WHEN x"81" => state_after_sub(I) <= x"0c";
					WHEN x"82" => state_after_sub(I) <= x"13";
					WHEN x"83" => state_after_sub(I) <= x"ec";
					WHEN x"84" => state_after_sub(I) <= x"5f";
					WHEN x"85" => state_after_sub(I) <= x"97";
					WHEN x"86" => state_after_sub(I) <= x"44";
					WHEN x"87" => state_after_sub(I) <= x"17";
					WHEN x"88" => state_after_sub(I) <= x"c4";
					WHEN x"89" => state_after_sub(I) <= x"a7";
					WHEN x"8a" => state_after_sub(I) <= x"7e";
					WHEN x"8b" => state_after_sub(I) <= x"3d";
					WHEN x"8c" => state_after_sub(I) <= x"64";
					WHEN x"8d" => state_after_sub(I) <= x"5d";
					WHEN x"8e" => state_after_sub(I) <= x"19";
					WHEN x"8f" => state_after_sub(I) <= x"73";  
					WHEN x"90" => state_after_sub(I) <= x"60";
					WHEN x"91" => state_after_sub(I) <= x"81";
					WHEN x"92" => state_after_sub(I) <= x"4f";
					WHEN x"93" => state_after_sub(I) <= x"dc";
					WHEN x"94" => state_after_sub(I) <= x"22";
					WHEN x"95" => state_after_sub(I) <= x"2a";
					WHEN x"96" => state_after_sub(I) <= x"90";
					WHEN x"97" => state_after_sub(I) <= x"88";
					WHEN x"98" => state_after_sub(I) <= x"46";
					WHEN x"99" => state_after_sub(I) <= x"ee";
					WHEN x"9a" => state_after_sub(I) <= x"b8";
					WHEN x"9b" => state_after_sub(I) <= x"14";
					WHEN x"9c" => state_after_sub(I) <= x"de";
					WHEN x"9d" => state_after_sub(I) <= x"5e";
					WHEN x"9e" => state_after_sub(I) <= x"0b";
					WHEN x"9f" => state_after_sub(I) <= x"db"; 
					WHEN x"a0" => state_after_sub(I) <= x"e0";
					WHEN x"a1" => state_after_sub(I) <= x"32";
					WHEN x"a2" => state_after_sub(I) <= x"3a";
					WHEN x"a3" => state_after_sub(I) <= x"0a";
					WHEN x"a4" => state_after_sub(I) <= x"49";
					WHEN x"a5" => state_after_sub(I) <= x"06";
					WHEN x"a6" => state_after_sub(I) <= x"24";
					WHEN x"a7" => state_after_sub(I) <= x"5c";
					WHEN x"a8" => state_after_sub(I) <= x"c2";
					WHEN x"a9" => state_after_sub(I) <= x"d3";
					WHEN x"aa" => state_after_sub(I) <= x"ac";
					WHEN x"ab" => state_after_sub(I) <= x"62";
					WHEN x"ac" => state_after_sub(I) <= x"91";
					WHEN x"ad" => state_after_sub(I) <= x"95";
					WHEN x"ae" => state_after_sub(I) <= x"e4";
					WHEN x"af" => state_after_sub(I) <= x"79";  
					WHEN x"b0" => state_after_sub(I) <= x"e7";
					WHEN x"b1" => state_after_sub(I) <= x"c8";
					WHEN x"b2" => state_after_sub(I) <= x"37";
					WHEN x"b3" => state_after_sub(I) <= x"6d";
					WHEN x"b4" => state_after_sub(I) <= x"8d";
					WHEN x"b5" => state_after_sub(I) <= x"d5";
					WHEN x"b6" => state_after_sub(I) <= x"4e";
					WHEN x"b7" => state_after_sub(I) <= x"a9";
					WHEN x"b8" => state_after_sub(I) <= x"6c";
					WHEN x"b9" => state_after_sub(I) <= x"56";
					WHEN x"ba" => state_after_sub(I) <= x"f4";
					WHEN x"bb" => state_after_sub(I) <= x"ea";
					WHEN x"bc" => state_after_sub(I) <= x"65";
					WHEN x"bd" => state_after_sub(I) <= x"7a";
					WHEN x"be" => state_after_sub(I) <= x"ae";
					WHEN x"bf" => state_after_sub(I) <= x"08";
					WHEN x"c0" => state_after_sub(I) <= x"ba";
					WHEN x"c1" => state_after_sub(I) <= x"78";
					WHEN x"c2" => state_after_sub(I) <= x"25";
					WHEN x"c3" => state_after_sub(I) <= x"2e";
					WHEN x"c4" => state_after_sub(I) <= x"1c";
					WHEN x"c5" => state_after_sub(I) <= x"a6";
					WHEN x"c6" => state_after_sub(I) <= x"b4";
					WHEN x"c7" => state_after_sub(I) <= x"c6";
					WHEN x"c8" => state_after_sub(I) <= x"e8";
					WHEN x"c9" => state_after_sub(I) <= x"dd";
					WHEN x"ca" => state_after_sub(I) <= x"74";
					WHEN x"cb" => state_after_sub(I) <= x"1f";
					WHEN x"cc" => state_after_sub(I) <= x"4b";
					WHEN x"cd" => state_after_sub(I) <= x"bd";
					WHEN x"ce" => state_after_sub(I) <= x"8b";
					WHEN x"cf" => state_after_sub(I) <= x"8a";  
					WHEN x"d0" => state_after_sub(I) <= x"70";
					WHEN x"d1" => state_after_sub(I) <= x"3e";
					WHEN x"d2" => state_after_sub(I) <= x"b5";
					WHEN x"d3" => state_after_sub(I) <= x"66";
					WHEN x"d4" => state_after_sub(I) <= x"48";
					WHEN x"d5" => state_after_sub(I) <= x"03";
					WHEN x"d6" => state_after_sub(I) <= x"f6";
					WHEN x"d7" => state_after_sub(I) <= x"0e";
					WHEN x"d8" => state_after_sub(I) <= x"61";
					WHEN x"d9" => state_after_sub(I) <= x"35";
					WHEN x"da" => state_after_sub(I) <= x"57";
					WHEN x"db" => state_after_sub(I) <= x"b9";
					WHEN x"dc" => state_after_sub(I) <= x"86";
					WHEN x"dd" => state_after_sub(I) <= x"c1";
					WHEN x"de" => state_after_sub(I) <= x"1d";
					WHEN x"df" => state_after_sub(I) <= x"9e"; 
					WHEN x"e0" => state_after_sub(I) <= x"e1";
					WHEN x"e1" => state_after_sub(I) <= x"f8";
					WHEN x"e2" => state_after_sub(I) <= x"98";
					WHEN x"e3" => state_after_sub(I) <= x"11";
					WHEN x"e4" => state_after_sub(I) <= x"69";
					WHEN x"e5" => state_after_sub(I) <= x"d9";
					WHEN x"e6" => state_after_sub(I) <= x"8e";
					WHEN x"e7" => state_after_sub(I) <= x"94";
					WHEN x"e8" => state_after_sub(I) <= x"9b";
					WHEN x"e9" => state_after_sub(I) <= x"1e";
					WHEN x"ea" => state_after_sub(I) <= x"87";
					WHEN x"eb" => state_after_sub(I) <= x"e9";
					WHEN x"ec" => state_after_sub(I) <= x"ce";
					WHEN x"ed" => state_after_sub(I) <= x"55";
					WHEN x"ee" => state_after_sub(I) <= x"28";
					WHEN x"ef" => state_after_sub(I) <= x"df";  
					WHEN x"f0" => state_after_sub(I) <= x"8c";
					WHEN x"f1" => state_after_sub(I) <= x"a1";
					WHEN x"f2" => state_after_sub(I) <= x"89";
					WHEN x"f3" => state_after_sub(I) <= x"0d";
					WHEN x"f4" => state_after_sub(I) <= x"bf";
					WHEN x"f5" => state_after_sub(I) <= x"e6";
					WHEN x"f6" => state_after_sub(I) <= x"42";
					WHEN x"f7" => state_after_sub(I) <= x"68";
					WHEN x"f8" => state_after_sub(I) <= x"41";
					WHEN x"f9" => state_after_sub(I) <= x"99";
					WHEN x"fa" => state_after_sub(I) <= x"2d";
					WHEN x"fb" => state_after_sub(I) <= x"0f";
					WHEN x"fc" => state_after_sub(I) <= x"b0";
					WHEN x"fd" => state_after_sub(I) <= x"54";
					WHEN x"fe" => state_after_sub(I) <= x"bb";
					WHEN x"ff" => state_after_sub(I) <= x"16";  
					WHEN others => null;  
				END CASE;   

	    --cWord <= state(I);
	    END LOOP;
  END PROCESS find;
--  state_after_sub <= t;
END rtl;
